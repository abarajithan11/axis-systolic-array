`timescale 1ns/1ps
`include "config.svh"

module top_ram_tb;
  localparam
    // Defined in config.svh
    R                   = `R                 ,
    C                   = `C                 ,
    WK                  = `WK                ,
    WX                  = `WX                ,
    WY                  = `WY                ,
    AXIL_BASE_ADDR      = `AXIL_BASE_ADDR    ,
    VALID_PROB          = `VALID_PROB        ,
    READY_PROB          = `READY_PROB        ,
    CLK_PERIOD          = `CLK_PERIOD        ,
    AXI_WIDTH           = `AXI_WIDTH         ,
    ADDR_WIDTH          = `ADDR_WIDTH        ,
    AXIL_WIDTH          = `AXIL_WIDTH        ,
    DIR                 = `DIR               ,
    WA                  = 32                 ,
    LM                  = 1                  ,
    LA                  = 1                  ,
    AXI_ID_WIDTH        = 6                  ,
    AXI_STRB_WIDTH      = AXI_WIDTH/8        ,
    AXI_MAX_BURST_LEN   = 32                 ,
    STRB_WIDTH          = 4                  ,
    DATA_WR_WIDTH       = AXIL_WIDTH         ,
    DATA_RD_WIDTH       = AXIL_WIDTH         ,
    LSB                 = $clog2(AXI_WIDTH)-3;


  // SIGNALS
  logic [ADDR_WIDTH     -1:0] reg_wr_addr;
  logic [AXIL_WIDTH     -1:0] reg_wr_data;
  logic [STRB_WIDTH     -1:0] reg_wr_strb;
  logic                       reg_wr_en  ;
  logic [ADDR_WIDTH     -1:0] reg_rd_addr;
  logic                       reg_rd_en  ;
  logic [AXIL_WIDTH     -1:0] reg_rd_data;

  logic                       mm2s_0_rd_en  ;
  logic [ADDR_WIDTH    -1:0]  mm2s_0_rd_addr;
  logic [AXI_WIDTH-1:0]       mm2s_0_rd_data;
  logic                       mm2s_0_rd_wait;
  logic                       mm2s_0_rd_ack ;
  logic                       mm2s_1_rd_en  ;
  logic [ADDR_WIDTH    -1:0]  mm2s_1_rd_addr;
  logic [AXI_WIDTH-1:0]       mm2s_1_rd_data;
  logic                       mm2s_1_rd_wait;
  logic                       mm2s_1_rd_ack ;
  logic                       mm2s_2_rd_en  ;
  logic [ADDR_WIDTH    -1:0]  mm2s_2_rd_addr;
  logic [AXI_WIDTH-1:0]       mm2s_2_rd_data;
  logic                       mm2s_2_rd_wait;
  logic                       mm2s_2_rd_ack ;
  logic                       s2mm_wr_en    ;
  logic [ADDR_WIDTH    -1:0]  s2mm_wr_addr  ;
  logic [AXI_WIDTH-1:0]       s2mm_wr_data  ;
  logic [AXI_STRB_WIDTH-1:0]  s2mm_wr_strb  ;
  logic                       s2mm_wr_wait  ;
  logic                       s2mm_wr_ack   ;

  top_sa_ram #(
    .R                 (R                ), 
    .C                 (C                ), 
    .WK                (WK               ), 
    .WX                (WX               ), 
    .WA                (WA               ), 
    .WY                (WY               ), 
    .LM                (LM               ), 
    .LA                (LA               ), 
    .AXI_WIDTH         (AXI_WIDTH        ), 
    .AXI_ID_WIDTH      (AXI_ID_WIDTH     ), 
    .AXI_STRB_WIDTH    (AXI_STRB_WIDTH   ), 
    .AXI_MAX_BURST_LEN (AXI_MAX_BURST_LEN), 
    .ADDR_WIDTH        (ADDR_WIDTH       ), 
    .AXIL_WIDTH        (AXIL_WIDTH       ), 
    .STRB_WIDTH        (STRB_WIDTH       ), 
    .AXIL_BASE_ADDR    (AXIL_BASE_ADDR   ) 
  ) dut(.*);

  logic clk = 0, rstn;
  initial forever #(CLK_PERIOD/2) clk = ~clk;

`ifdef VERILATOR
  `define AUTOMATIC
`else
  `define AUTOMATIC automatic
`endif

  export "DPI-C" task _get_config;
  export "DPI-C" task set_config;
  import "DPI-C" context task get_byte_a32 (input int unsigned addr, output byte data);
  import "DPI-C" context task set_byte_a32 (input int unsigned addr, input byte data);
  import "DPI-C" context function chandle get_mp ();
  import "DPI-C" context task `AUTOMATIC run(input chandle mem_ptr_virtual, input chandle p_config, ref int done);
  // import "DPI-C" context task void print_output (chandle mem_ptr_virtual);


  task automatic _get_config(input chandle config_base, input int offset, output int data);
    data = dut.CONTROLLER.cfg [offset];
  endtask

  task automatic set_config(input chandle config_base, input int offset, input int data);
    dut.CONTROLLER.cfg [offset] <= data;
  endtask

  int done = 0;
  byte tmp_byte_0, tmp_byte_1, tmp_byte_2;

  always_comb begin
    mm2s_0_rd_wait = 0;
    mm2s_0_rd_ack  = 1;
    mm2s_0_rd_data = '0;
    tmp_byte_0     = 0;
    if (mm2s_0_rd_en) begin
      for (int i = 0; i < AXI_WIDTH/8; i++) begin
        get_byte_a32((mm2s_0_rd_addr) + i, tmp_byte_0);
        mm2s_0_rd_data[i*8 +: 8] = tmp_byte_0;
      end
    end

    mm2s_1_rd_wait = 0;
    mm2s_1_rd_ack  = 1;
    mm2s_1_rd_data = '0;
    tmp_byte_1     = 0;
    if (mm2s_1_rd_en) begin
      for (int i = 0; i < AXI_WIDTH/8; i++) begin
        get_byte_a32((mm2s_1_rd_addr) + i, tmp_byte_1);
        mm2s_1_rd_data[i*8 +: 8] = tmp_byte_1;
      end
    end

    mm2s_2_rd_wait = 0;
    mm2s_2_rd_ack  = 1;
    mm2s_2_rd_data = '0;
    tmp_byte_2     = 0;
    if (mm2s_2_rd_en) begin
      for (int i = 0; i < AXI_WIDTH/8; i++) begin
        get_byte_a32((32'(mm2s_2_rd_addr)) + i, tmp_byte_2);
        mm2s_2_rd_data[i*8 +: 8] = tmp_byte_2;
      end
    end
  end

  always_ff @(posedge clk) begin : Axi_rw
    s2mm_wr_wait <= 0;
    s2mm_wr_ack  <= s2mm_wr_en;
    if (s2mm_wr_en) 
      for (int i = 0; i < AXI_WIDTH/8; i++) 
        if (s2mm_wr_strb[i]) 
          set_byte_a32((32'(s2mm_wr_addr)) + i, s2mm_wr_data[i*8 +: 8]);
  end
  
  initial begin
    $dumpfile("top_tb.vcd");
    $dumpvars();
    #1000us;
    $fatal(1, "\n\nError: Timeout \n\n");
  end

  int file_out, file_exp, status, error=0, i=0;
  byte out_byte, exp_byte;

  chandle mem_ptr_virtual, cfg_ptr_virtual;
  initial begin
    rstn <= 0;
    repeat(2) @(posedge clk) #10ps;
    rstn <= 1;
    mem_ptr_virtual = get_mp();
    
    while (done == 0) begin
      run(mem_ptr_virtual, cfg_ptr_virtual, done);
      @(posedge clk) #10ps;
    end
    done = 0;


    // Read from output & expected and compare
    file_out = $fopen({DIR, "/y.bin"}, "rb");
    file_exp = $fopen({DIR, "/y_exp.bin" }, "rb");
    if (file_out==0 || file_exp==0) $fatal(0, "Error: Failed to open output/expected file(s).");

    while($feof(file_exp) == 0) begin
      if ($feof(file_out)) $fatal(0, "Error: output file is shorter than expected file.");
      else begin
        out_byte = $fgetc(file_out);
        exp_byte = $fgetc(file_exp);
        // Compare
        if (exp_byte != out_byte) begin
          $display("Mismatch at index %0d: Expected %h, Found %h", i, exp_byte, out_byte);
          error += 1;
        end 
      end
      i += 1;
    end
    $fclose(file_exp);
    $fclose(file_out);
    
    if (error==0) $display("\n\nVerification successful: Output matches Expected data. \nError count: %0d\n\n", error);
    else          $fatal (0, "\n\nERROR: Output data does not match Expected data.\n\n");
    $finish;
  end

endmodule
